// ---------------------------
// 1. Behavioral Modeling
// ---------------------------
module full_adder_behavioral(
    input a, b, cin,
    output reg sum, cout
);
    always @(*) begin
        {cout, sum} = a + b + cin;  
    end
endmodule

// ---------------------------
// 2. Dataflow (RTL) Modeling
// ---------------------------
module full_adder_dataflow(
    input a, b, cin,
    output sum, cout
);
    assign sum  = a ^ b ^ cin;                        
    assign cout = (a & b) | (b & cin) | (a & cin);    
endmodule

// ---------------------------
// 3. Structural Modeling
// ---------------------------
module full_adder_structural(
    input a, b, cin,
    output sum, cout
);
    wire w1, w2, w3;

    // Half Adder 1
    xor (w1, a, b);        
    and (w2, a, b);        

    // Half Adder 2
    xor (sum, w1, cin);    
    and (w3, w1, cin);     

    // Final carry
    or (cout, w2, w3);
endmodule
